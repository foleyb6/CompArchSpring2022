module RAM(Addr, RW, DataI, DataO);

input [31:0] Addr;
input RW;
input [31:0] DataI;
output reg [31:0] DataO;

reg [31:0] RAM0, RAM1, RAM2, RAM3, RAM4, RAM5, RAM6, RAM7, RAM8, RAM9;
reg [31:0] RAM10, RAM11, RAM12, RAM13, RAM14, RAM15, RAM16, RAM17, RAM18, RAM19;
reg [31:0] RAM20, RAM21, RAM22, RAM23, RAM24, RAM25, RAM26, RAM27, RAM28, RAM29;
reg [31:0] RAM30, RAM31, RAM32, RAM33, RAM34, RAM35, RAM36, RAM37, RAM38, RAM39;
reg [31:0] RAM40, RAM41, RAM42, RAM43, RAM44, RAM45, RAM46, RAM47, RAM48, RAM49;
reg [31:0] RAM50, RAM51, RAM52, RAM53, RAM54, RAM55, RAM56, RAM57, RAM58, RAM59;
reg [31:0] RAM60, RAM61, RAM62, RAM63, RAM64, RAM65, RAM66, RAM67, RAM68, RAM69;
reg [31:0] RAM70, RAM71, RAM72, RAM73, RAM74, RAM75, RAM76, RAM77, RAM78, RAM79;
reg [31:0] RAM80, RAM81, RAM82, RAM83, RAM84, RAM85, RAM86, RAM87, RAM88, RAM89;
reg [31:0] RAM90, RAM91, RAM92, RAM93, RAM94, RAM95, RAM96, RAM97, RAM98, RAM99;
reg [31:0] RAM100, RAM101, RAM102, RAM103, RAM104, RAM105, RAM106, RAM107, RAM108, RAM109;
reg [31:0] RAM110, RAM111, RAM112, RAM113, RAM114, RAM115, RAM116, RAM117, RAM118, RAM119;
reg [31:0] RAM120, RAM121, RAM122, RAM123, RAM124, RAM125, RAM126, RAM127, RAM128, RAM129;
reg [31:0] RAM130, RAM131, RAM132, RAM133, RAM134, RAM135, RAM136, RAM137, RAM138, RAM139;
reg [31:0] RAM140, RAM141, RAM142, RAM143, RAM144, RAM145, RAM146, RAM147, RAM148, RAM149;
reg [31:0] RAM150, RAM151, RAM152, RAM153, RAM154, RAM155, RAM156, RAM157, RAM158, RAM159;
reg [31:0] RAM160, RAM161, RAM162, RAM163, RAM164, RAM165, RAM166, RAM167, RAM168, RAM169;
reg [31:0] RAM170, RAM171, RAM172, RAM173, RAM174, RAM175, RAM176, RAM177, RAM178, RAM179;
reg [31:0] RAM180, RAM181, RAM182, RAM183, RAM184, RAM185, RAM186, RAM187, RAM188, RAM189;
reg [31:0] RAM190, RAM191, RAM192, RAM193, RAM194, RAM195, RAM196, RAM197, RAM198, RAM199;
reg [31:0] RAM200, RAM201, RAM202, RAM203, RAM204, RAM205, RAM206, RAM207, RAM208, RAM209;
reg [31:0] RAM210, RAM211, RAM212, RAM213, RAM214, RAM215, RAM216, RAM217, RAM218, RAM219;
reg [31:0] RAM220, RAM221, RAM222, RAM223, RAM224, RAM225, RAM226, RAM227, RAM228, RAM229;
reg [31:0] RAM230, RAM231, RAM232, RAM233, RAM234, RAM235, RAM236, RAM237, RAM238, RAM239;
reg [31:0] RAM240, RAM241, RAM242, RAM243, RAM244, RAM245, RAM246, RAM247, RAM248, RAM249;
reg [31:0] RAM250, RAM251, RAM252, RAM253, RAM254, RAM255;

always @(RW)
begin
	case(Addr)
	32'd0 : RAM0 <= DataI;
	32'd1 : RAM1 <= DataI;
	32'd2 : RAM2 <= DataI;
	32'd3 : RAM3 <= DataI;
	32'd4 : RAM4 <= DataI;
	32'd5 : RAM5 <= DataI;
	32'd6 : RAM6 <= DataI;
	32'd7 : RAM7 <= DataI;
	32'd8 : RAM8 <= DataI;
	32'd9 : RAM9 <= DataI;
	32'd10 : RAM10 <= DataI;
	32'd11 : RAM11 <= DataI;
	32'd12 : RAM12 <= DataI;
	32'd13 : RAM13 <= DataI;
	32'd14 : RAM14 <= DataI;
	32'd15 : RAM15 <= DataI;
	32'd16 : RAM16 <= DataI;
	32'd17 : RAM17 <= DataI;
	32'd18 : RAM18 <= DataI;
	32'd19 : RAM19 <= DataI;
	32'd20 : RAM20 <= DataI;
	32'd21 : RAM21 <= DataI;
	32'd22 : RAM22 <= DataI;
	32'd23 : RAM23 <= DataI;
	32'd24 : RAM24 <= DataI;
	32'd25 : RAM25 <= DataI;
	32'd26 : RAM26 <= DataI;
	32'd27 : RAM27 <= DataI;
	32'd28 : RAM28 <= DataI;
	32'd29 : RAM29 <= DataI;
	32'd30 : RAM30 <= DataI;
	32'd31 : RAM31 <= DataI;
	32'd32 : RAM32 <= DataI;
	32'd33 : RAM33 <= DataI;
	32'd34 : RAM34 <= DataI;
	32'd35 : RAM35 <= DataI;
	32'd36 : RAM36 <= DataI;
	32'd37 : RAM37 <= DataI;
	32'd38 : RAM38 <= DataI;
	32'd39 : RAM39 <= DataI;
	32'd40 : RAM40 <= DataI;
	32'd41 : RAM41 <= DataI;
	32'd42 : RAM42 <= DataI;
	32'd43 : RAM43 <= DataI;
	32'd44 : RAM44 <= DataI;
	32'd45 : RAM45 <= DataI;
	32'd46 : RAM46 <= DataI;
	32'd47 : RAM47 <= DataI;
	32'd48 : RAM48 <= DataI;
	32'd49 : RAM49 <= DataI;
	32'd50 : RAM50 <= DataI;
	32'd51 : RAM51 <= DataI;
	32'd52 : RAM52 <= DataI;
	32'd53 : RAM53 <= DataI;
	32'd54 : RAM54 <= DataI;
	32'd55 : RAM55 <= DataI;
	32'd56 : RAM56 <= DataI;
	32'd57 : RAM57 <= DataI;
	32'd58 : RAM58 <= DataI;
	32'd59 : RAM59 <= DataI;
	32'd60 : RAM60 <= DataI;
	32'd61 : RAM61 <= DataI;
	32'd62 : RAM62 <= DataI;
	32'd63 : RAM63 <= DataI;
	32'd64 : RAM64 <= DataI;
	32'd65 : RAM65 <= DataI;
	32'd66 : RAM66 <= DataI;
	32'd67 : RAM67 <= DataI;
	32'd68 : RAM68 <= DataI;
	32'd69 : RAM69 <= DataI;
	32'd70 : RAM70 <= DataI;
	32'd71 : RAM71 <= DataI;
	32'd72 : RAM72 <= DataI;
	32'd73 : RAM73 <= DataI;
	32'd74 : RAM74 <= DataI;
	32'd75 : RAM75 <= DataI;
	32'd76 : RAM76 <= DataI;
	32'd77 : RAM77 <= DataI;
	32'd78 : RAM78 <= DataI;
	32'd79 : RAM79 <= DataI;
	32'd80 : RAM80 <= DataI;
	32'd81 : RAM81 <= DataI;
	32'd82 : RAM82 <= DataI;
	32'd83 : RAM83 <= DataI;
	32'd84 : RAM84 <= DataI;
	32'd85 : RAM85 <= DataI;
	32'd86 : RAM86 <= DataI;
	32'd87 : RAM87 <= DataI;
	32'd88 : RAM88 <= DataI;
	32'd89 : RAM89 <= DataI;
	32'd90 : RAM90 <= DataI;
	32'd91 : RAM91 <= DataI;
	32'd92 : RAM92 <= DataI;
	32'd93 : RAM93 <= DataI;
	32'd94 : RAM94 <= DataI;
	32'd95 : RAM95 <= DataI;
	32'd96 : RAM96 <= DataI;
	32'd97 : RAM97 <= DataI;
	32'd98 : RAM98 <= DataI;
	32'd99 : RAM99 <= DataI;
	32'd100 : RAM100 <= DataI;
	32'd101 : RAM101 <= DataI;
	32'd102 : RAM102 <= DataI;
	32'd103 : RAM103 <= DataI;
	32'd104 : RAM104 <= DataI;
	32'd105 : RAM105 <= DataI;
	32'd106 : RAM106 <= DataI;
	32'd107 : RAM107 <= DataI;
	32'd108 : RAM108 <= DataI;
	32'd109 : RAM109 <= DataI;
	32'd110 : RAM110 <= DataI;
	32'd111 : RAM111 <= DataI;
	32'd112 : RAM112 <= DataI;
	32'd113 : RAM113 <= DataI;
	32'd114 : RAM114 <= DataI;
	32'd115 : RAM115 <= DataI;
	32'd116 : RAM116 <= DataI;
	32'd117 : RAM117 <= DataI;
	32'd118 : RAM118 <= DataI;
	32'd119 : RAM119 <= DataI;
	32'd120 : RAM120 <= DataI;
	32'd121 : RAM121 <= DataI;
	32'd122 : RAM122 <= DataI;
	32'd123 : RAM123 <= DataI;
	32'd124 : RAM124 <= DataI;
	32'd125 : RAM125 <= DataI;
	32'd126 : RAM126 <= DataI;
	32'd127 : RAM127 <= DataI;
	32'd128 : RAM128 <= DataI;
	32'd129 : RAM129 <= DataI;
	32'd130 : RAM130 <= DataI;
	32'd131 : RAM131 <= DataI;
	32'd132 : RAM132 <= DataI;
	32'd133 : RAM133 <= DataI;
	32'd134 : RAM134 <= DataI;
	32'd135 : RAM135 <= DataI;
	32'd136 : RAM136 <= DataI;
	32'd137 : RAM137 <= DataI;
	32'd138 : RAM138 <= DataI;
	32'd139 : RAM139 <= DataI;
	32'd140 : RAM140 <= DataI;
	32'd141 : RAM141 <= DataI;
	32'd142 : RAM142 <= DataI;
	32'd143 : RAM143 <= DataI;
	32'd144 : RAM144 <= DataI;
	32'd145 : RAM145 <= DataI;
	32'd146 : RAM146 <= DataI;
	32'd147 : RAM147 <= DataI;
	32'd148 : RAM148 <= DataI;
	32'd149 : RAM149 <= DataI;
	32'd150 : RAM150 <= DataI;
	32'd151 : RAM151 <= DataI;
	32'd152 : RAM152 <= DataI;
	32'd153 : RAM153 <= DataI;
	32'd154 : RAM154 <= DataI;
	32'd155 : RAM155 <= DataI;
	32'd156 : RAM156 <= DataI;
	32'd157 : RAM157 <= DataI;
	32'd158 : RAM158 <= DataI;
	32'd159 : RAM159 <= DataI;
	32'd160 : RAM160 <= DataI;
	32'd161 : RAM161 <= DataI;
	32'd162 : RAM162 <= DataI;
	32'd163 : RAM163 <= DataI;
	32'd164 : RAM164 <= DataI;
	32'd165 : RAM165 <= DataI;
	32'd166 : RAM166 <= DataI;
	32'd167 : RAM167 <= DataI;
	32'd168 : RAM168 <= DataI;
	32'd169 : RAM169 <= DataI;
	32'd170 : RAM170 <= DataI;
	32'd171 : RAM171 <= DataI;
	32'd172 : RAM172 <= DataI;
	32'd173 : RAM173 <= DataI;
	32'd174 : RAM174 <= DataI;
	32'd175 : RAM175 <= DataI;
	32'd176 : RAM176 <= DataI;
	32'd177 : RAM177 <= DataI;
	32'd178 : RAM178 <= DataI;
	32'd179 : RAM179 <= DataI;
	32'd180 : RAM180 <= DataI;
	32'd181 : RAM181 <= DataI;
	32'd182 : RAM182 <= DataI;
	32'd183 : RAM183 <= DataI;
	32'd184 : RAM184 <= DataI;
	32'd185 : RAM185 <= DataI;
	32'd186 : RAM186 <= DataI;
	32'd187 : RAM187 <= DataI;
	32'd188 : RAM188 <= DataI;
	32'd189 : RAM189 <= DataI;
	32'd190 : RAM190 <= DataI;
	32'd191 : RAM191 <= DataI;
	32'd192 : RAM192 <= DataI;
	32'd193 : RAM193 <= DataI;
	32'd194 : RAM194 <= DataI;
	32'd195 : RAM195 <= DataI;
	32'd196 : RAM196 <= DataI;
	32'd197 : RAM197 <= DataI;
	32'd198 : RAM198 <= DataI;
	32'd199 : RAM199 <= DataI;
	32'd200 : RAM200 <= DataI;
	32'd201 : RAM201 <= DataI;
	32'd202 : RAM202 <= DataI;
	32'd203 : RAM203 <= DataI;
	32'd204 : RAM204 <= DataI;
	32'd205 : RAM205 <= DataI;
	32'd206 : RAM206 <= DataI;
	32'd207 : RAM207 <= DataI;
	32'd208 : RAM208 <= DataI;
	32'd209 : RAM209 <= DataI;
	32'd210 : RAM210 <= DataI;
	32'd211 : RAM211 <= DataI;
	32'd212 : RAM212 <= DataI;
	32'd213 : RAM213 <= DataI;
	32'd214 : RAM214 <= DataI;
	32'd215 : RAM215 <= DataI;
	32'd216 : RAM216 <= DataI;
	32'd217 : RAM217 <= DataI;
	32'd218 : RAM218 <= DataI;
	32'd219 : RAM219 <= DataI;
	32'd220 : RAM220 <= DataI;
	32'd221 : RAM221 <= DataI;
	32'd222 : RAM222 <= DataI;
	32'd223 : RAM223 <= DataI;
	32'd224 : RAM224 <= DataI;
	32'd225 : RAM225 <= DataI;
	32'd226 : RAM226 <= DataI;
	32'd227 : RAM227 <= DataI;
	32'd228 : RAM228 <= DataI;
	32'd229 : RAM229 <= DataI;
	32'd230 : RAM230 <= DataI;
	32'd231 : RAM231 <= DataI;
	32'd232 : RAM232 <= DataI;
	32'd233 : RAM233 <= DataI;
	32'd234 : RAM234 <= DataI;
	32'd235 : RAM235 <= DataI;
	32'd236 : RAM236 <= DataI;
	32'd237 : RAM237 <= DataI;
	32'd238 : RAM238 <= DataI;
	32'd239 : RAM239 <= DataI;
	32'd240 : RAM240 <= DataI;
	32'd241 : RAM241 <= DataI;
	32'd242 : RAM242 <= DataI;
	32'd243 : RAM243 <= DataI;
	32'd244 : RAM244 <= DataI;
	32'd245 : RAM245 <= DataI;
	32'd246 : RAM246 <= DataI;
	32'd247 : RAM247 <= DataI;
	32'd248 : RAM248 <= DataI;
	32'd249 : RAM249 <= DataI;
	32'd250 : RAM250 <= DataI;
	32'd251 : RAM251 <= DataI;
	32'd252 : RAM252 <= DataI;
	32'd253 : RAM253 <= DataI;
	32'd254 : RAM254 <= DataI;
	32'd255 : RAM255 <= DataI;
	endcase
end

always @(RW)
begin
	case(Addr)
	32'd0:DataO <= RAM0;
	32'd1:DataO <= RAM1;
	32'd2:DataO <= RAM2;
	32'd3:DataO <= RAM3;
	32'd4:DataO <= RAM4;
	32'd5:DataO <= RAM5;
	32'd6:DataO <= RAM6;
	32'd7:DataO <= RAM7;
	32'd8:DataO <= RAM8;
	32'd9:DataO <= RAM9;
	32'd10:DataO <= RAM10;
	32'd11:DataO <= RAM11;
	32'd12:DataO <= RAM12;
	32'd13:DataO <= RAM13;
	32'd14:DataO <= RAM14;
	32'd15:DataO <= RAM15;
	32'd16:DataO <= RAM16;
	32'd17:DataO <= RAM17;
	32'd18:DataO <= RAM18;
	32'd19:DataO <= RAM19;
	32'd20:DataO <= RAM20;
	32'd21:DataO <= RAM21;
	32'd22:DataO <= RAM22;
	32'd23:DataO <= RAM23;
	32'd24:DataO <= RAM24;
	32'd25:DataO <= RAM25;
	32'd26:DataO <= RAM26;
	32'd27:DataO <= RAM27;
	32'd28:DataO <= RAM28;
	32'd29:DataO <= RAM29;
	32'd30:DataO <= RAM30;
	32'd31:DataO <= RAM31;
	32'd32:DataO <= RAM32;
	32'd33:DataO <= RAM33;
	32'd34:DataO <= RAM34;
	32'd35:DataO <= RAM35;
	32'd36:DataO <= RAM36;
	32'd37:DataO <= RAM37;
	32'd38:DataO <= RAM38;
	32'd39:DataO <= RAM39;
	32'd40:DataO <= RAM40;
	32'd41:DataO <= RAM41;
	32'd42:DataO <= RAM42;
	32'd43:DataO <= RAM43;
	32'd44:DataO <= RAM44;
	32'd45:DataO <= RAM45;
	32'd46:DataO <= RAM46;
	32'd47:DataO <= RAM47;
	32'd48:DataO <= RAM48;
	32'd49:DataO <= RAM49;
	32'd50:DataO <= RAM50;
	32'd51:DataO <= RAM51;
	32'd52:DataO <= RAM52;
	32'd53:DataO <= RAM53;
	32'd54:DataO <= RAM54;
	32'd55:DataO <= RAM55;
	32'd56:DataO <= RAM56;
	32'd57:DataO <= RAM57;
	32'd58:DataO <= RAM58;
	32'd59:DataO <= RAM59;
	32'd60:DataO <= RAM60;
	32'd61:DataO <= RAM61;
	32'd62:DataO <= RAM62;
	32'd63:DataO <= RAM63;
	32'd64:DataO <= RAM64;
	32'd65:DataO <= RAM65;
	32'd66:DataO <= RAM66;
	32'd67:DataO <= RAM67;
	32'd68:DataO <= RAM68;
	32'd69:DataO <= RAM69;
	32'd70:DataO <= RAM70;
	32'd71:DataO <= RAM71;
	32'd72:DataO <= RAM72;
	32'd73:DataO <= RAM73;
	32'd74:DataO <= RAM74;
	32'd75:DataO <= RAM75;
	32'd76:DataO <= RAM76;
	32'd77:DataO <= RAM77;
	32'd78:DataO <= RAM78;
	32'd79:DataO <= RAM79;
	32'd80:DataO <= RAM80;
	32'd81:DataO <= RAM81;
	32'd82:DataO <= RAM82;
	32'd83:DataO <= RAM83;
	32'd84:DataO <= RAM84;
	32'd85:DataO <= RAM85;
	32'd86:DataO <= RAM86;
	32'd87:DataO <= RAM87;
	32'd88:DataO <= RAM88;
	32'd89:DataO <= RAM89;
	32'd90:DataO <= RAM90;
	32'd91:DataO <= RAM91;
	32'd92:DataO <= RAM92;
	32'd93:DataO <= RAM93;
	32'd94:DataO <= RAM94;
	32'd95:DataO <= RAM95;
	32'd96:DataO <= RAM96;
	32'd97:DataO <= RAM97;
	32'd98:DataO <= RAM98;
	32'd99:DataO <= RAM99;
	32'd100:DataO <= RAM100;
	32'd101:DataO <= RAM101;
	32'd102:DataO <= RAM102;
	32'd103:DataO <= RAM103;
	32'd104:DataO <= RAM104;
	32'd105:DataO <= RAM105;
	32'd106:DataO <= RAM106;
	32'd107:DataO <= RAM107;
	32'd108:DataO <= RAM108;
	32'd109:DataO <= RAM109;
	32'd110:DataO <= RAM110;
	32'd111:DataO <= RAM111;
	32'd112:DataO <= RAM112;
	32'd113:DataO <= RAM113;
	32'd114:DataO <= RAM114;
	32'd115:DataO <= RAM115;
	32'd116:DataO <= RAM116;
	32'd117:DataO <= RAM117;
	32'd118:DataO <= RAM118;
	32'd119:DataO <= RAM119;
	32'd120:DataO <= RAM120;
	32'd121:DataO <= RAM121;
	32'd122:DataO <= RAM122;
	32'd123:DataO <= RAM123;
	32'd124:DataO <= RAM124;
	32'd125:DataO <= RAM125;
	32'd126:DataO <= RAM126;
	32'd127:DataO <= RAM127;
	32'd128:DataO <= RAM128;
	32'd129:DataO <= RAM129;
	32'd130:DataO <= RAM130;
	32'd131:DataO <= RAM131;
	32'd132:DataO <= RAM132;
	32'd133:DataO <= RAM133;
	32'd134:DataO <= RAM134;
	32'd135:DataO <= RAM135;
	32'd136:DataO <= RAM136;
	32'd137:DataO <= RAM137;
	32'd138:DataO <= RAM138;
	32'd139:DataO <= RAM139;
	32'd140:DataO <= RAM140;
	32'd141:DataO <= RAM141;
	32'd142:DataO <= RAM142;
	32'd143:DataO <= RAM143;
	32'd144:DataO <= RAM144;
	32'd145:DataO <= RAM145;
	32'd146:DataO <= RAM146;
	32'd147:DataO <= RAM147;
	32'd148:DataO <= RAM148;
	32'd149:DataO <= RAM149;
	32'd150:DataO <= RAM150;
	32'd151:DataO <= RAM151;
	32'd152:DataO <= RAM152;
	32'd153:DataO <= RAM153;
	32'd154:DataO <= RAM154;
	32'd155:DataO <= RAM155;
	32'd156:DataO <= RAM156;
	32'd157:DataO <= RAM157;
	32'd158:DataO <= RAM158;
	32'd159:DataO <= RAM159;
	32'd160:DataO <= RAM160;
	32'd161:DataO <= RAM161;
	32'd162:DataO <= RAM162;
	32'd163:DataO <= RAM163;
	32'd164:DataO <= RAM164;
	32'd165:DataO <= RAM165;
	32'd166:DataO <= RAM166;
	32'd167:DataO <= RAM167;
	32'd168:DataO <= RAM168;
	32'd169:DataO <= RAM169;
	32'd170:DataO <= RAM170;
	32'd171:DataO <= RAM171;
	32'd172:DataO <= RAM172;
	32'd173:DataO <= RAM173;
	32'd174:DataO <= RAM174;
	32'd175:DataO <= RAM175;
	32'd176:DataO <= RAM176;
	32'd177:DataO <= RAM177;
	32'd178:DataO <= RAM178;
	32'd179:DataO <= RAM179;
	32'd180:DataO <= RAM180;
	32'd181:DataO <= RAM181;
	32'd182:DataO <= RAM182;
	32'd183:DataO <= RAM183;
	32'd184:DataO <= RAM184;
	32'd185:DataO <= RAM185;
	32'd186:DataO <= RAM186;
	32'd187:DataO <= RAM187;
	32'd188:DataO <= RAM188;
	32'd189:DataO <= RAM189;
	32'd190:DataO <= RAM190;
	32'd191:DataO <= RAM191;
	32'd192:DataO <= RAM192;
	32'd193:DataO <= RAM193;
	32'd194:DataO <= RAM194;
	32'd195:DataO <= RAM195;
	32'd196:DataO <= RAM196;
	32'd197:DataO <= RAM197;
	32'd198:DataO <= RAM198;
	32'd199:DataO <= RAM199;
	32'd200:DataO <= RAM200;
	32'd201:DataO <= RAM201;
	32'd202:DataO <= RAM202;
	32'd203:DataO <= RAM203;
	32'd204:DataO <= RAM204;
	32'd205:DataO <= RAM205;
	32'd206:DataO <= RAM206;
	32'd207:DataO <= RAM207;
	32'd208:DataO <= RAM208;
	32'd209:DataO <= RAM209;
	32'd210:DataO <= RAM210;
	32'd211:DataO <= RAM211;
	32'd212:DataO <= RAM212;
	32'd213:DataO <= RAM213;
	32'd214:DataO <= RAM214;
	32'd215:DataO <= RAM215;
	32'd216:DataO <= RAM216;
	32'd217:DataO <= RAM217;
	32'd218:DataO <= RAM218;
	32'd219:DataO <= RAM219;
	32'd220:DataO <= RAM220;
	32'd221:DataO <= RAM221;
	32'd222:DataO <= RAM222;
	32'd223:DataO <= RAM223;
	32'd224:DataO <= RAM224;
	32'd225:DataO <= RAM225;
	32'd226:DataO <= RAM226;
	32'd227:DataO <= RAM227;
	32'd228:DataO <= RAM228;
	32'd229:DataO <= RAM229;
	32'd230:DataO <= RAM230;
	32'd231:DataO <= RAM231;
	32'd232:DataO <= RAM232;
	32'd233:DataO <= RAM233;
	32'd234:DataO <= RAM234;
	32'd235:DataO <= RAM235;
	32'd236:DataO <= RAM236;
	32'd237:DataO <= RAM237;
	32'd238:DataO <= RAM238;
	32'd239:DataO <= RAM239;
	32'd240:DataO <= RAM240;
	32'd241:DataO <= RAM241;
	32'd242:DataO <= RAM242;
	32'd243:DataO <= RAM243;
	32'd244:DataO <= RAM244;
	32'd245:DataO <= RAM245;
	32'd246:DataO <= RAM246;
	32'd247:DataO <= RAM247;
	32'd248:DataO <= RAM248;
	32'd249:DataO <= RAM249;
	32'd250:DataO <= RAM250;
	32'd251:DataO <= RAM251;
	32'd252:DataO <= RAM252;
	32'd253:DataO <= RAM253;
	32'd254:DataO <= RAM254;
	32'd255:DataO <= RAM255;
	endcase
end

endmodule
