module RAM(Addr, RAMW, RAMR, Input, Output);

input [31:0] Addr;
input RAMW, RAMR;
input [31:0] Input;
output reg [31:0] Output;

reg [31:0] RAM0, RAM1, RAM2, RAM3, RAM4, RAM5, RAM6, RAM7, RAM8, RAM9;
reg [31:0] RAM10, RAM11, RAM12, RAM13, RAM14, RAM15, RAM16, RAM17, RAM18, RAM19;
reg [31:0] RAM20, RAM21, RAM22, RAM23, RAM24, RAM25, RAM26, RAM27, RAM28, RAM29;
reg [31:0] RAM30, RAM31, RAM32, RAM33, RAM34, RAM35, RAM36, RAM37, RAM38, RAM39;
reg [31:0] RAM40, RAM41, RAM42, RAM43, RAM44, RAM45, RAM46, RAM47, RAM48, RAM49;
reg [31:0] RAM50, RAM51, RAM52, RAM53, RAM54, RAM55, RAM56, RAM57, RAM58, RAM59;
reg [31:0] RAM60, RAM61, RAM62, RAM63, RAM64, RAM65, RAM66, RAM67, RAM68, RAM69;
reg [31:0] RAM70, RAM71, RAM72, RAM73, RAM74, RAM75, RAM76, RAM77, RAM78, RAM79;
reg [31:0] RAM80, RAM81, RAM82, RAM83, RAM84, RAM85, RAM86, RAM87, RAM88, RAM89;
reg [31:0] RAM90, RAM91, RAM92, RAM93, RAM94, RAM95, RAM96, RAM97, RAM98, RAM99;
reg [31:0] RAM100, RAM101, RAM102, RAM103, RAM104, RAM105, RAM106, RAM107, RAM108, RAM109;
reg [31:0] RAM110, RAM111, RAM112, RAM113, RAM114, RAM115, RAM116, RAM117, RAM118, RAM119;
reg [31:0] RAM120, RAM121, RAM122, RAM123, RAM124, RAM125, RAM126, RAM127, RAM128, RAM129;
reg [31:0] RAM130, RAM131, RAM132, RAM133, RAM134, RAM135, RAM136, RAM137, RAM138, RAM139;
reg [31:0] RAM140, RAM141, RAM142, RAM143, RAM144, RAM145, RAM146, RAM147, RAM148, RAM149;
reg [31:0] RAM150, RAM151, RAM152, RAM153, RAM154, RAM155, RAM156, RAM157, RAM158, RAM159;
reg [31:0] RAM160, RAM161, RAM162, RAM163, RAM164, RAM165, RAM166, RAM167, RAM168, RAM169;
reg [31:0] RAM170, RAM171, RAM172, RAM173, RAM174, RAM175, RAM176, RAM177, RAM178, RAM179;
reg [31:0] RAM180, RAM181, RAM182, RAM183, RAM184, RAM185, RAM186, RAM187, RAM188, RAM189;
reg [31:0] RAM190, RAM191, RAM192, RAM193, RAM194, RAM195, RAM196, RAM197, RAM198, RAM199;
reg [31:0] RAM200, RAM201, RAM202, RAM203, RAM204, RAM205, RAM206, RAM207, RAM208, RAM209;
reg [31:0] RAM210, RAM211, RAM212, RAM213, RAM214, RAM215, RAM216, RAM217, RAM218, RAM219;
reg [31:0] RAM220, RAM221, RAM222, RAM223, RAM224, RAM225, RAM226, RAM227, RAM228, RAM229;
reg [31:0] RAM230, RAM231, RAM232, RAM233, RAM234, RAM235, RAM236, RAM237, RAM238, RAM239;
reg [31:0] RAM240, RAM241, RAM242, RAM243, RAM244, RAM245, RAM246, RAM247, RAM248, RAM249;
reg [31:0] RAM250, RAM251, RAM252, RAM253, RAM254, RAM255;

always @(RAMW)
begin
	case(Addr)
	32'd0 : RAM0 <= Input;
	32'd1 : RAM1 <= Input;
	32'd2 : RAM2 <= Input;
	32'd3 : RAM3 <= Input;
	32'd4 : RAM4 <= Input;
	32'd5 : RAM5 <= Input;
	32'd6 : RAM6 <= Input;
	32'd7 : RAM7 <= Input;
	32'd8 : RAM8 <= Input;
	32'd9 : RAM9 <= Input;
	32'd10 : RAM10 <= Input;
	32'd11 : RAM11 <= Input;
	32'd12 : RAM12 <= Input;
	32'd13 : RAM13 <= Input;
	32'd14 : RAM14 <= Input;
	32'd15 : RAM15 <= Input;
	32'd16 : RAM16 <= Input;
	32'd17 : RAM17 <= Input;
	32'd18 : RAM18 <= Input;
	32'd19 : RAM19 <= Input;
	32'd20 : RAM20 <= Input;
	32'd21 : RAM21 <= Input;
	32'd22 : RAM22 <= Input;
	32'd23 : RAM23 <= Input;
	32'd24 : RAM24 <= Input;
	32'd25 : RAM25 <= Input;
	32'd26 : RAM26 <= Input;
	32'd27 : RAM27 <= Input;
	32'd28 : RAM28 <= Input;
	32'd29 : RAM29 <= Input;
	32'd30 : RAM30 <= Input;
	32'd31 : RAM31 <= Input;
	32'd32 : RAM32 <= Input;
	32'd33 : RAM33 <= Input;
	32'd34 : RAM34 <= Input;
	32'd35 : RAM35 <= Input;
	32'd36 : RAM36 <= Input;
	32'd37 : RAM37 <= Input;
	32'd38 : RAM38 <= Input;
	32'd39 : RAM39 <= Input;
	32'd40 : RAM40 <= Input;
	32'd41 : RAM41 <= Input;
	32'd42 : RAM42 <= Input;
	32'd43 : RAM43 <= Input;
	32'd44 : RAM44 <= Input;
	32'd45 : RAM45 <= Input;
	32'd46 : RAM46 <= Input;
	32'd47 : RAM47 <= Input;
	32'd48 : RAM48 <= Input;
	32'd49 : RAM49 <= Input;
	32'd50 : RAM50 <= Input;
	32'd51 : RAM51 <= Input;
	32'd52 : RAM52 <= Input;
	32'd53 : RAM53 <= Input;
	32'd54 : RAM54 <= Input;
	32'd55 : RAM55 <= Input;
	32'd56 : RAM56 <= Input;
	32'd57 : RAM57 <= Input;
	32'd58 : RAM58 <= Input;
	32'd59 : RAM59 <= Input;
	32'd60 : RAM60 <= Input;
	32'd61 : RAM61 <= Input;
	32'd62 : RAM62 <= Input;
	32'd63 : RAM63 <= Input;
	32'd64 : RAM64 <= Input;
	32'd65 : RAM65 <= Input;
	32'd66 : RAM66 <= Input;
	32'd67 : RAM67 <= Input;
	32'd68 : RAM68 <= Input;
	32'd69 : RAM69 <= Input;
	32'd70 : RAM70 <= Input;
	32'd71 : RAM71 <= Input;
	32'd72 : RAM72 <= Input;
	32'd73 : RAM73 <= Input;
	32'd74 : RAM74 <= Input;
	32'd75 : RAM75 <= Input;
	32'd76 : RAM76 <= Input;
	32'd77 : RAM77 <= Input;
	32'd78 : RAM78 <= Input;
	32'd79 : RAM79 <= Input;
	32'd80 : RAM80 <= Input;
	32'd81 : RAM81 <= Input;
	32'd82 : RAM82 <= Input;
	32'd83 : RAM83 <= Input;
	32'd84 : RAM84 <= Input;
	32'd85 : RAM85 <= Input;
	32'd86 : RAM86 <= Input;
	32'd87 : RAM87 <= Input;
	32'd88 : RAM88 <= Input;
	32'd89 : RAM89 <= Input;
	32'd90 : RAM90 <= Input;
	32'd91 : RAM91 <= Input;
	32'd92 : RAM92 <= Input;
	32'd93 : RAM93 <= Input;
	32'd94 : RAM94 <= Input;
	32'd95 : RAM95 <= Input;
	32'd96 : RAM96 <= Input;
	32'd97 : RAM97 <= Input;
	32'd98 : RAM98 <= Input;
	32'd99 : RAM99 <= Input;
	32'd100 : RAM100 <= Input;
	32'd101 : RAM101 <= Input;
	32'd102 : RAM102 <= Input;
	32'd103 : RAM103 <= Input;
	32'd104 : RAM104 <= Input;
	32'd105 : RAM105 <= Input;
	32'd106 : RAM106 <= Input;
	32'd107 : RAM107 <= Input;
	32'd108 : RAM108 <= Input;
	32'd109 : RAM109 <= Input;
	32'd110 : RAM110 <= Input;
	32'd111 : RAM111 <= Input;
	32'd112 : RAM112 <= Input;
	32'd113 : RAM113 <= Input;
	32'd114 : RAM114 <= Input;
	32'd115 : RAM115 <= Input;
	32'd116 : RAM116 <= Input;
	32'd117 : RAM117 <= Input;
	32'd118 : RAM118 <= Input;
	32'd119 : RAM119 <= Input;
	32'd120 : RAM120 <= Input;
	32'd121 : RAM121 <= Input;
	32'd122 : RAM122 <= Input;
	32'd123 : RAM123 <= Input;
	32'd124 : RAM124 <= Input;
	32'd125 : RAM125 <= Input;
	32'd126 : RAM126 <= Input;
	32'd127 : RAM127 <= Input;
	32'd128 : RAM128 <= Input;
	32'd129 : RAM129 <= Input;
	32'd130 : RAM130 <= Input;
	32'd131 : RAM131 <= Input;
	32'd132 : RAM132 <= Input;
	32'd133 : RAM133 <= Input;
	32'd134 : RAM134 <= Input;
	32'd135 : RAM135 <= Input;
	32'd136 : RAM136 <= Input;
	32'd137 : RAM137 <= Input;
	32'd138 : RAM138 <= Input;
	32'd139 : RAM139 <= Input;
	32'd140 : RAM140 <= Input;
	32'd141 : RAM141 <= Input;
	32'd142 : RAM142 <= Input;
	32'd143 : RAM143 <= Input;
	32'd144 : RAM144 <= Input;
	32'd145 : RAM145 <= Input;
	32'd146 : RAM146 <= Input;
	32'd147 : RAM147 <= Input;
	32'd148 : RAM148 <= Input;
	32'd149 : RAM149 <= Input;
	32'd150 : RAM150 <= Input;
	32'd151 : RAM151 <= Input;
	32'd152 : RAM152 <= Input;
	32'd153 : RAM153 <= Input;
	32'd154 : RAM154 <= Input;
	32'd155 : RAM155 <= Input;
	32'd156 : RAM156 <= Input;
	32'd157 : RAM157 <= Input;
	32'd158 : RAM158 <= Input;
	32'd159 : RAM159 <= Input;
	32'd160 : RAM160 <= Input;
	32'd161 : RAM161 <= Input;
	32'd162 : RAM162 <= Input;
	32'd163 : RAM163 <= Input;
	32'd164 : RAM164 <= Input;
	32'd165 : RAM165 <= Input;
	32'd166 : RAM166 <= Input;
	32'd167 : RAM167 <= Input;
	32'd168 : RAM168 <= Input;
	32'd169 : RAM169 <= Input;
	32'd170 : RAM170 <= Input;
	32'd171 : RAM171 <= Input;
	32'd172 : RAM172 <= Input;
	32'd173 : RAM173 <= Input;
	32'd174 : RAM174 <= Input;
	32'd175 : RAM175 <= Input;
	32'd176 : RAM176 <= Input;
	32'd177 : RAM177 <= Input;
	32'd178 : RAM178 <= Input;
	32'd179 : RAM179 <= Input;
	32'd180 : RAM180 <= Input;
	32'd181 : RAM181 <= Input;
	32'd182 : RAM182 <= Input;
	32'd183 : RAM183 <= Input;
	32'd184 : RAM184 <= Input;
	32'd185 : RAM185 <= Input;
	32'd186 : RAM186 <= Input;
	32'd187 : RAM187 <= Input;
	32'd188 : RAM188 <= Input;
	32'd189 : RAM189 <= Input;
	32'd190 : RAM190 <= Input;
	32'd191 : RAM191 <= Input;
	32'd192 : RAM192 <= Input;
	32'd193 : RAM193 <= Input;
	32'd194 : RAM194 <= Input;
	32'd195 : RAM195 <= Input;
	32'd196 : RAM196 <= Input;
	32'd197 : RAM197 <= Input;
	32'd198 : RAM198 <= Input;
	32'd199 : RAM199 <= Input;
	32'd200 : RAM200 <= Input;
	32'd201 : RAM201 <= Input;
	32'd202 : RAM202 <= Input;
	32'd203 : RAM203 <= Input;
	32'd204 : RAM204 <= Input;
	32'd205 : RAM205 <= Input;
	32'd206 : RAM206 <= Input;
	32'd207 : RAM207 <= Input;
	32'd208 : RAM208 <= Input;
	32'd209 : RAM209 <= Input;
	32'd210 : RAM210 <= Input;
	32'd211 : RAM211 <= Input;
	32'd212 : RAM212 <= Input;
	32'd213 : RAM213 <= Input;
	32'd214 : RAM214 <= Input;
	32'd215 : RAM215 <= Input;
	32'd216 : RAM216 <= Input;
	32'd217 : RAM217 <= Input;
	32'd218 : RAM218 <= Input;
	32'd219 : RAM219 <= Input;
	32'd220 : RAM220 <= Input;
	32'd221 : RAM221 <= Input;
	32'd222 : RAM222 <= Input;
	32'd223 : RAM223 <= Input;
	32'd224 : RAM224 <= Input;
	32'd225 : RAM225 <= Input;
	32'd226 : RAM226 <= Input;
	32'd227 : RAM227 <= Input;
	32'd228 : RAM228 <= Input;
	32'd229 : RAM229 <= Input;
	32'd230 : RAM230 <= Input;
	32'd231 : RAM231 <= Input;
	32'd232 : RAM232 <= Input;
	32'd233 : RAM233 <= Input;
	32'd234 : RAM234 <= Input;
	32'd235 : RAM235 <= Input;
	32'd236 : RAM236 <= Input;
	32'd237 : RAM237 <= Input;
	32'd238 : RAM238 <= Input;
	32'd239 : RAM239 <= Input;
	32'd240 : RAM240 <= Input;
	32'd241 : RAM241 <= Input;
	32'd242 : RAM242 <= Input;
	32'd243 : RAM243 <= Input;
	32'd244 : RAM244 <= Input;
	32'd245 : RAM245 <= Input;
	32'd246 : RAM246 <= Input;
	32'd247 : RAM247 <= Input;
	32'd248 : RAM248 <= Input;
	32'd249 : RAM249 <= Input;
	32'd250 : RAM250 <= Input;
	32'd251 : RAM251 <= Input;
	32'd252 : RAM252 <= Input;
	32'd253 : RAM253 <= Input;
	32'd254 : RAM254 <= Input;
	32'd255 : RAM255 <= Input;
	endcase
end

always @(RAMR)
begin
	case(Addr)
	32'd0:Output <= RAM0;
	32'd1:Output <= RAM1;
	32'd2:Output <= RAM2;
	32'd3:Output <= RAM3;
	32'd4:Output <= RAM4;
	32'd5:Output <= RAM5;
	32'd6:Output <= RAM6;
	32'd7:Output <= RAM7;
	32'd8:Output <= RAM8;
	32'd9:Output <= RAM9;
	32'd10:Output <= RAM10;
	32'd11:Output <= RAM11;
	32'd12:Output <= RAM12;
	32'd13:Output <= RAM13;
	32'd14:Output <= RAM14;
	32'd15:Output <= RAM15;
	32'd16:Output <= RAM16;
	32'd17:Output <= RAM17;
	32'd18:Output <= RAM18;
	32'd19:Output <= RAM19;
	32'd20:Output <= RAM20;
	32'd21:Output <= RAM21;
	32'd22:Output <= RAM22;
	32'd23:Output <= RAM23;
	32'd24:Output <= RAM24;
	32'd25:Output <= RAM25;
	32'd26:Output <= RAM26;
	32'd27:Output <= RAM27;
	32'd28:Output <= RAM28;
	32'd29:Output <= RAM29;
	32'd30:Output <= RAM30;
	32'd31:Output <= RAM31;
	32'd32:Output <= RAM32;
	32'd33:Output <= RAM33;
	32'd34:Output <= RAM34;
	32'd35:Output <= RAM35;
	32'd36:Output <= RAM36;
	32'd37:Output <= RAM37;
	32'd38:Output <= RAM38;
	32'd39:Output <= RAM39;
	32'd40:Output <= RAM40;
	32'd41:Output <= RAM41;
	32'd42:Output <= RAM42;
	32'd43:Output <= RAM43;
	32'd44:Output <= RAM44;
	32'd45:Output <= RAM45;
	32'd46:Output <= RAM46;
	32'd47:Output <= RAM47;
	32'd48:Output <= RAM48;
	32'd49:Output <= RAM49;
	32'd50:Output <= RAM50;
	32'd51:Output <= RAM51;
	32'd52:Output <= RAM52;
	32'd53:Output <= RAM53;
	32'd54:Output <= RAM54;
	32'd55:Output <= RAM55;
	32'd56:Output <= RAM56;
	32'd57:Output <= RAM57;
	32'd58:Output <= RAM58;
	32'd59:Output <= RAM59;
	32'd60:Output <= RAM60;
	32'd61:Output <= RAM61;
	32'd62:Output <= RAM62;
	32'd63:Output <= RAM63;
	32'd64:Output <= RAM64;
	32'd65:Output <= RAM65;
	32'd66:Output <= RAM66;
	32'd67:Output <= RAM67;
	32'd68:Output <= RAM68;
	32'd69:Output <= RAM69;
	32'd70:Output <= RAM70;
	32'd71:Output <= RAM71;
	32'd72:Output <= RAM72;
	32'd73:Output <= RAM73;
	32'd74:Output <= RAM74;
	32'd75:Output <= RAM75;
	32'd76:Output <= RAM76;
	32'd77:Output <= RAM77;
	32'd78:Output <= RAM78;
	32'd79:Output <= RAM79;
	32'd80:Output <= RAM80;
	32'd81:Output <= RAM81;
	32'd82:Output <= RAM82;
	32'd83:Output <= RAM83;
	32'd84:Output <= RAM84;
	32'd85:Output <= RAM85;
	32'd86:Output <= RAM86;
	32'd87:Output <= RAM87;
	32'd88:Output <= RAM88;
	32'd89:Output <= RAM89;
	32'd90:Output <= RAM90;
	32'd91:Output <= RAM91;
	32'd92:Output <= RAM92;
	32'd93:Output <= RAM93;
	32'd94:Output <= RAM94;
	32'd95:Output <= RAM95;
	32'd96:Output <= RAM96;
	32'd97:Output <= RAM97;
	32'd98:Output <= RAM98;
	32'd99:Output <= RAM99;
	32'd100:Output <= RAM100;
	32'd101:Output <= RAM101;
	32'd102:Output <= RAM102;
	32'd103:Output <= RAM103;
	32'd104:Output <= RAM104;
	32'd105:Output <= RAM105;
	32'd106:Output <= RAM106;
	32'd107:Output <= RAM107;
	32'd108:Output <= RAM108;
	32'd109:Output <= RAM109;
	32'd110:Output <= RAM110;
	32'd111:Output <= RAM111;
	32'd112:Output <= RAM112;
	32'd113:Output <= RAM113;
	32'd114:Output <= RAM114;
	32'd115:Output <= RAM115;
	32'd116:Output <= RAM116;
	32'd117:Output <= RAM117;
	32'd118:Output <= RAM118;
	32'd119:Output <= RAM119;
	32'd120:Output <= RAM120;
	32'd121:Output <= RAM121;
	32'd122:Output <= RAM122;
	32'd123:Output <= RAM123;
	32'd124:Output <= RAM124;
	32'd125:Output <= RAM125;
	32'd126:Output <= RAM126;
	32'd127:Output <= RAM127;
	32'd128:Output <= RAM128;
	32'd129:Output <= RAM129;
	32'd130:Output <= RAM130;
	32'd131:Output <= RAM131;
	32'd132:Output <= RAM132;
	32'd133:Output <= RAM133;
	32'd134:Output <= RAM134;
	32'd135:Output <= RAM135;
	32'd136:Output <= RAM136;
	32'd137:Output <= RAM137;
	32'd138:Output <= RAM138;
	32'd139:Output <= RAM139;
	32'd140:Output <= RAM140;
	32'd141:Output <= RAM141;
	32'd142:Output <= RAM142;
	32'd143:Output <= RAM143;
	32'd144:Output <= RAM144;
	32'd145:Output <= RAM145;
	32'd146:Output <= RAM146;
	32'd147:Output <= RAM147;
	32'd148:Output <= RAM148;
	32'd149:Output <= RAM149;
	32'd150:Output <= RAM150;
	32'd151:Output <= RAM151;
	32'd152:Output <= RAM152;
	32'd153:Output <= RAM153;
	32'd154:Output <= RAM154;
	32'd155:Output <= RAM155;
	32'd156:Output <= RAM156;
	32'd157:Output <= RAM157;
	32'd158:Output <= RAM158;
	32'd159:Output <= RAM159;
	32'd160:Output <= RAM160;
	32'd161:Output <= RAM161;
	32'd162:Output <= RAM162;
	32'd163:Output <= RAM163;
	32'd164:Output <= RAM164;
	32'd165:Output <= RAM165;
	32'd166:Output <= RAM166;
	32'd167:Output <= RAM167;
	32'd168:Output <= RAM168;
	32'd169:Output <= RAM169;
	32'd170:Output <= RAM170;
	32'd171:Output <= RAM171;
	32'd172:Output <= RAM172;
	32'd173:Output <= RAM173;
	32'd174:Output <= RAM174;
	32'd175:Output <= RAM175;
	32'd176:Output <= RAM176;
	32'd177:Output <= RAM177;
	32'd178:Output <= RAM178;
	32'd179:Output <= RAM179;
	32'd180:Output <= RAM180;
	32'd181:Output <= RAM181;
	32'd182:Output <= RAM182;
	32'd183:Output <= RAM183;
	32'd184:Output <= RAM184;
	32'd185:Output <= RAM185;
	32'd186:Output <= RAM186;
	32'd187:Output <= RAM187;
	32'd188:Output <= RAM188;
	32'd189:Output <= RAM189;
	32'd190:Output <= RAM190;
	32'd191:Output <= RAM191;
	32'd192:Output <= RAM192;
	32'd193:Output <= RAM193;
	32'd194:Output <= RAM194;
	32'd195:Output <= RAM195;
	32'd196:Output <= RAM196;
	32'd197:Output <= RAM197;
	32'd198:Output <= RAM198;
	32'd199:Output <= RAM199;
	32'd200:Output <= RAM200;
	32'd201:Output <= RAM201;
	32'd202:Output <= RAM202;
	32'd203:Output <= RAM203;
	32'd204:Output <= RAM204;
	32'd205:Output <= RAM205;
	32'd206:Output <= RAM206;
	32'd207:Output <= RAM207;
	32'd208:Output <= RAM208;
	32'd209:Output <= RAM209;
	32'd210:Output <= RAM210;
	32'd211:Output <= RAM211;
	32'd212:Output <= RAM212;
	32'd213:Output <= RAM213;
	32'd214:Output <= RAM214;
	32'd215:Output <= RAM215;
	32'd216:Output <= RAM216;
	32'd217:Output <= RAM217;
	32'd218:Output <= RAM218;
	32'd219:Output <= RAM219;
	32'd220:Output <= RAM220;
	32'd221:Output <= RAM221;
	32'd222:Output <= RAM222;
	32'd223:Output <= RAM223;
	32'd224:Output <= RAM224;
	32'd225:Output <= RAM225;
	32'd226:Output <= RAM226;
	32'd227:Output <= RAM227;
	32'd228:Output <= RAM228;
	32'd229:Output <= RAM229;
	32'd230:Output <= RAM230;
	32'd231:Output <= RAM231;
	32'd232:Output <= RAM232;
	32'd233:Output <= RAM233;
	32'd234:Output <= RAM234;
	32'd235:Output <= RAM235;
	32'd236:Output <= RAM236;
	32'd237:Output <= RAM237;
	32'd238:Output <= RAM238;
	32'd239:Output <= RAM239;
	32'd240:Output <= RAM240;
	32'd241:Output <= RAM241;
	32'd242:Output <= RAM242;
	32'd243:Output <= RAM243;
	32'd244:Output <= RAM244;
	32'd245:Output <= RAM245;
	32'd246:Output <= RAM246;
	32'd247:Output <= RAM247;
	32'd248:Output <= RAM248;
	32'd249:Output <= RAM249;
	32'd250:Output <= RAM250;
	32'd251:Output <= RAM251;
	32'd252:Output <= RAM252;
	32'd253:Output <= RAM253;
	32'd254:Output <= RAM254;
	32'd255:Output <= RAM255;
	endcase
end

endmodule
