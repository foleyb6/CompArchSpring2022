module Decoder(Selector, WriAdd, WriEn, Clock);
input [4:0] WriAdd;
input WriEn, Clock;

output reg [31:0] Selector;


always @(posedge Clock)
if(WriEn == 1)
begin
	case(WriAdd)
	5'b00000 : Selector = 32'b00000000000000000000000000000001;
	5'b00001 : Selector = 32'b00000000000000000000000000000010;
	5'b00010 : Selector = 32'b00000000000000000000000000000100;
	5'b00011 : Selector = 32'b00000000000000000000000000001000;
	5'b00100 : Selector = 32'b00000000000000000000000000010000;
	5'b00101 : Selector = 32'b00000000000000000000000000100000;
	5'b00110 : Selector = 32'b00000000000000000000000001000000;
	5'b00111 : Selector = 32'b00000000000000000000000010000000;
	5'b01000 : Selector = 32'b00000000000000000000000100000000;
	5'b01001 : Selector = 32'b00000000000000000000001000000000;
	5'b01010 : Selector = 32'b00000000000000000000010000000000;
	5'b01011 : Selector = 32'b00000000000000000000100000000000;
	5'b01100 : Selector = 32'b00000000000000000001000000000000;
	5'b01101 : Selector = 32'b00000000000000000010000000000000;
	5'b01110 : Selector = 32'b00000000000000000100000000000000;
	5'b01111 : Selector = 32'b00000000000000001000000000000000;
	5'b10000 : Selector = 32'b00000000000000010000000000000000;
	5'b10001 : Selector = 32'b00000000000000100000000000000000;
	5'b10010 : Selector = 32'b00000000000001000000000000000000;
	5'b10011 : Selector = 32'b00000000000010000000000000000000;
	5'b10100 : Selector = 32'b00000000000100000000000000000000;
	5'b10101 : Selector = 32'b00000000001000000000000000000000;
	5'b10110 : Selector = 32'b00000000010000000000000000000000;
	5'b10111 : Selector = 32'b00000000100000000000000000000000;
	5'b11000 : Selector = 32'b00000001000000000000000000000000;
	5'b11001 : Selector = 32'b00000010000000000000000000000000;
	5'b11010 : Selector = 32'b00000100000000000000000000000000;
	5'b11011 : Selector = 32'b00001000000000000000000000000000;
	5'b11100 : Selector = 32'b00010000000000000000000000000000;
	5'b11101 : Selector = 32'b00100000000000000000000000000000;
	5'b11110 : Selector = 32'b01000000000000000000000000000000;
	5'b11111 : Selector = 32'b10000000000000000000000000000000;
	endcase
end
else
begin
Selector = 32'b00000000000000000000000000000000;
end

endmodule
